------------------------------------------
-----------COMANDOS PARA LCD--------------
------------�NO MODIFICAR!---------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

package COMANDOS_LCD_REVB is

FUNCTION LCD_INI(DATO : STD_LOGIC_VECTOR(1 DOWNTO 0)) RETURN STD_LOGIC_VECTOR;
FUNCTION CHAR(DATO1 : STRING) RETURN STD_LOGIC_VECTOR;
FUNCTION POS(DATO2,DATO3 : INTEGER) RETURN STD_LOGIC_VECTOR;
FUNCTION CD_SHIFT(DATO4,DATO5 : INTEGER) RETURN STD_LOGIC_VECTOR;
FUNCTION CHAR_ASCII(DATO6 : STD_LOGIC_VECTOR(7 DOWNTO 0))RETURN STD_LOGIC_VECTOR;
FUNCTION CODIGO_FIN(DATO7 : INTEGER) RETURN STD_LOGIC_VECTOR;
FUNCTION BUCLE_INI(DATO8 : INTEGER)RETURN STD_LOGIC_VECTOR;
FUNCTION BUCLE_FIN(DATO9 : INTEGER)RETURN STD_LOGIC_VECTOR;
FUNCTION INT_NUM(DATO10 : INTEGER)RETURN STD_LOGIC_VECTOR;
---
FUNCTION CREAR_CHAR(DATO11: INTEGER)RETURN STD_LOGIC_VECTOR;--DATAOUT8

FUNCTION CHAR_CREADO(DATO12: INTEGER)RETURN STD_LOGIC_VECTOR;--DATAOUT9

FUNCTION LIMPIAR_PANTALLA(DATO9 : STD_LOGIC)RETURN STD_LOGIC_VECTOR;

CONSTANT a:STRING:="a";CONSTANT j:STRING:="j";CONSTANT s:STRING:="s";
CONSTANT b:STRING:="b";CONSTANT k:STRING:="k";CONSTANT t:STRING:="t";
CONSTANT c:STRING:="c";CONSTANT l:STRING:="l";CONSTANT u:STRING:="u";
CONSTANT d:STRING:="d";CONSTANT m:STRING:="m";CONSTANT v:STRING:="v";
CONSTANT e:STRING:="e";CONSTANT n:STRING:="n";CONSTANT w:STRING:="w";
CONSTANT f:STRING:="f";CONSTANT o:STRING:="o";CONSTANT x:STRING:="x";
CONSTANT g:STRING:="g";CONSTANT p:STRING:="p";CONSTANT y:STRING:="y";
CONSTANT h:STRING:="h";CONSTANT q:STRING:="q";CONSTANT z:STRING:="z";
CONSTANT i:STRING:="i";CONSTANT r:STRING:="r";

CONSTANT Ma:STRING:="A";CONSTANT Mj:STRING:="J";CONSTANT MAs:STRING:="S";
CONSTANT Mb:STRING:="B";CONSTANT Mk:STRING:="K";CONSTANT Mt:STRING:="T";
CONSTANT Mc:STRING:="C";CONSTANT Ml:STRING:="L";CONSTANT Mu:STRING:="U";
CONSTANT Md:STRING:="D";CONSTANT Mm:STRING:="M";CONSTANT Mv:STRING:="V";
CONSTANT Me:STRING:="E";CONSTANT Mn:STRING:="N";CONSTANT Mw:STRING:="W";
CONSTANT Mf:STRING:="F";CONSTANT Mo:STRING:="O";CONSTANT Mx:STRING:="X";
CONSTANT Mg:STRING:="G";CONSTANT Mp:STRING:="P";CONSTANT My:STRING:="Y";
CONSTANT Mh:STRING:="H";CONSTANT Mq:STRING:="Q";CONSTANT Mz:STRING:="Z";
CONSTANT Mi:STRING:="I";CONSTANT Mr:STRING:="R";


CONSTANT N1:STRING:="1";CONSTANT N5:STRING:="5";CONSTANT N9:STRING:="9";
CONSTANT N2:STRING:="2";CONSTANT N6:STRING:="6";CONSTANT N0:STRING:="0";
CONSTANT N3:STRING:="3";CONSTANT N7:STRING:="7";
CONSTANT N4:STRING:="4";CONSTANT N8:STRING:="8";

end COMANDOS_LCD_REVB;

package body COMANDOS_LCD_REVB is

----LCD_INI()------
-------------------
FUNCTION LCD_INI(DATO : STD_LOGIC_VECTOR(1 DOWNTO 0)) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
CASE DATO IS
WHEN "00" => RETURN '1'&x"01";
WHEN "01" => RETURN '1'&x"02";
WHEN "10" => RETURN '1'&x"03";
WHEN OTHERS => RETURN '1'&x"04";
END CASE;
END LCD_INI;
-----------------

-----CHAR()-----
-----------------
FUNCTION CHAR(DATO1 : STRING) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT1 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
CASE DATO1 IS
WHEN a => RETURN '1'&x"09";
WHEN b => RETURN '1'&x"0A";
WHEN c => RETURN '1'&x"0B";
WHEN d => RETURN '1'&x"0C";
WHEN e => RETURN '1'&x"0D";
WHEN f => RETURN '1'&x"0E";
WHEN g => RETURN '1'&x"0F";
WHEN h => RETURN '1'&x"10";
WHEN i => RETURN '1'&x"11";
WHEN j => RETURN '1'&x"12";
WHEN k => RETURN '1'&x"13";
WHEN l => RETURN '1'&x"14";
WHEN m => RETURN '1'&x"15";
WHEN n => RETURN '1'&x"16";
WHEN o => RETURN '1'&x"17";
WHEN p => RETURN '1'&x"18";
WHEN q => RETURN '1'&x"19";
WHEN r => RETURN '1'&x"1A";
WHEN s => RETURN '1'&x"1B";
WHEN t => RETURN '1'&x"1C";
WHEN u => RETURN '1'&x"1D";
WHEN v => RETURN '1'&x"1E";
WHEN w => RETURN '1'&x"1F";
WHEN x => RETURN '1'&x"20";
WHEN y => RETURN '1'&x"21";
WHEN z => RETURN '1'&x"22";
----
WHEN MA => RETURN '1'&x"23";
WHEN MB => RETURN '1'&x"24";
WHEN MC => RETURN '1'&x"25";
WHEN MD => RETURN '1'&x"26";
WHEN ME => RETURN '1'&x"27";
WHEN MF => RETURN '1'&x"28";
WHEN MG => RETURN '1'&x"29";
WHEN MH => RETURN '1'&x"2A";
WHEN MI => RETURN '1'&x"2B";
WHEN MJ => RETURN '1'&x"2C";
WHEN MK => RETURN '1'&x"2D";
WHEN ML => RETURN '1'&x"2E";
WHEN MM => RETURN '1'&x"2F";
WHEN MN => RETURN '1'&x"30";
WHEN MO => RETURN '1'&x"31";
WHEN MP => RETURN '1'&x"32";
WHEN MQ => RETURN '1'&x"33";
WHEN MR => RETURN '1'&x"34";
WHEN MAS => RETURN '1'&x"35";
WHEN MT => RETURN '1'&x"36";
WHEN MU => RETURN '1'&x"37";
WHEN MV => RETURN '1'&x"38";
WHEN MW => RETURN '1'&x"39";
WHEN MX => RETURN '1'&x"3A";
WHEN MY => RETURN '1'&x"3B";
WHEN MZ => RETURN '1'&x"3C";
----
WHEN N0 => RETURN '1'&x"3D";
WHEN N1 => RETURN '1'&x"3E";
WHEN N2 => RETURN '1'&x"3F";
WHEN N3 => RETURN '1'&x"40";
WHEN N4 => RETURN '1'&x"41";
WHEN N5 => RETURN '1'&x"42";
WHEN N6 => RETURN '1'&x"43";
WHEN N7 => RETURN '1'&x"44";
WHEN N8 => RETURN '1'&x"45";
WHEN N9 => RETURN '1'&x"46";
WHEN OTHERS => RETURN '1'&x"47";
END CASE;
END CHAR;
  
---INT_NUM()----
----------------

FUNCTION INT_NUM(DATO10 : INTEGER) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT6 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
CASE DATO10 IS
WHEN 0 => RETURN '0'&x"30";
WHEN 1 => RETURN '0'&x"31";
WHEN 2 => RETURN '0'&x"32";
WHEN 3 => RETURN '0'&x"33";
WHEN 4 => RETURN '0'&x"34";
WHEN 5 => RETURN '0'&x"35";
WHEN 6 => RETURN '0'&x"36";
WHEN 7 => RETURN '0'&x"37";
WHEN 8 => RETURN '0'&x"38";
WHEN 9 => RETURN '0'&x"39";
WHEN OTHERS => RETURN '0'&x"30";
END CASE;
END INT_NUM;

----------------
  
----POS()------
--------------------
FUNCTION POS(DATO2,DATO3 : INTEGER) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT2 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF 	DATO2 = 1 AND DATO3 = 1  THEN RETURN '1'&x"50";
ELSIF DATO2 = 1 AND DATO3 = 2  THEN RETURN '1'&x"51";
ELSIF DATO2 = 1 AND DATO3 = 3  THEN RETURN '1'&x"52";
ELSIF DATO2 = 1 AND DATO3 = 4  THEN RETURN '1'&x"53";
ELSIF DATO2 = 1 AND DATO3 = 5  THEN RETURN '1'&x"54";
ELSIF DATO2 = 1 AND DATO3 = 6  THEN RETURN '1'&x"55";
ELSIF DATO2 = 1 AND DATO3 = 7  THEN RETURN '1'&x"56";
ELSIF DATO2 = 1 AND DATO3 = 8  THEN RETURN '1'&x"57";
ELSIF DATO2 = 1 AND DATO3 = 9  THEN RETURN '1'&x"58";
ELSIF DATO2 = 1 AND DATO3 = 10 THEN RETURN '1'&x"59";
ELSIF DATO2 = 1 AND DATO3 = 11 THEN RETURN '1'&x"5A";
ELSIF DATO2 = 1 AND DATO3 = 12 THEN RETURN '1'&x"5B";
ELSIF DATO2 = 1 AND DATO3 = 13 THEN RETURN '1'&x"5C";
ELSIF DATO2 = 1 AND DATO3 = 14 THEN RETURN '1'&x"5D";
ELSIF DATO2 = 1 AND DATO3 = 15 THEN RETURN '1'&x"5E";
ELSIF DATO2 = 1 AND DATO3 = 16 THEN RETURN '1'&x"5F";
ELSIF DATO2 = 1 AND DATO3 = 17 THEN RETURN '1'&x"60";
ELSIF DATO2 = 1 AND DATO3 = 18 THEN RETURN '1'&x"61";
ELSIF DATO2 = 1 AND DATO3 = 19 THEN RETURN '1'&x"62";
ELSIF DATO2 = 1 AND DATO3 = 20 THEN RETURN '1'&x"63";
-------
ELSIF	DATO2 = 2 AND DATO3 = 1  THEN RETURN '1'&x"64";
ELSIF DATO2 = 2 AND DATO3 = 2  THEN RETURN '1'&x"65";
ELSIF DATO2 = 2 AND DATO3 = 3  THEN RETURN '1'&x"66";
ELSIF DATO2 = 2 AND DATO3 = 4  THEN RETURN '1'&x"67";
ELSIF DATO2 = 2 AND DATO3 = 5  THEN RETURN '1'&x"68";
ELSIF DATO2 = 2 AND DATO3 = 6  THEN RETURN '1'&x"69";
ELSIF DATO2 = 2 AND DATO3 = 7  THEN RETURN '1'&x"6A";
ELSIF DATO2 = 2 AND DATO3 = 8  THEN RETURN '1'&x"6B";
ELSIF DATO2 = 2 AND DATO3 = 9  THEN RETURN '1'&x"6C";
ELSIF DATO2 = 2 AND DATO3 = 10 THEN RETURN '1'&x"6D";
ELSIF DATO2 = 2 AND DATO3 = 11 THEN RETURN '1'&x"6E";
ELSIF DATO2 = 2 AND DATO3 = 12 THEN RETURN '1'&x"6F";
ELSIF DATO2 = 2 AND DATO3 = 13 THEN RETURN '1'&x"70";
ELSIF DATO2 = 2 AND DATO3 = 14 THEN RETURN '1'&x"71";
ELSIF DATO2 = 2 AND DATO3 = 15 THEN RETURN '1'&x"72";
ELSIF DATO2 = 2 AND DATO3 = 16 THEN RETURN '1'&x"73";
ELSIF DATO2 = 2 AND DATO3 = 17 THEN RETURN '1'&x"74";
ELSIF DATO2 = 2 AND DATO3 = 18 THEN RETURN '1'&x"75";
ELSIF DATO2 = 2 AND DATO3 = 19 THEN RETURN '1'&x"76";
ELSIF DATO2 = 2 AND DATO3 = 20 THEN RETURN '1'&x"77";
ELSE RETURN '1'&x"77";
--ELSE NULL;
END IF;
END POS;
-------------------

----CD_SHIFT()------
--------------------
FUNCTION CD_SHIFT(DATO4,DATO5 : INTEGER) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT3 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF 	DATO4 = 0 AND DATO5 = 0  THEN RETURN '1'&x"78";
ELSIF DATO4 = 0 AND DATO5 = 1  THEN RETURN '1'&x"79";
ELSIF DATO4 = 1 AND DATO5 = 0  THEN RETURN '1'&x"7A";
ELSIF DATO4 = 1 AND DATO5 = 1  THEN RETURN '1'&x"7B";
--ELSE NULL;
ELSE RETURN '1'&x"7B";
END IF;
END CD_SHIFT;
-------------------

------BUCLE_INI()----
----------------------
FUNCTION BUCLE_INI(DATO8 : INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT6 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF DATO8 = 1 THEN RETURN '1'&x"7C";
ELSE RETURN '1'&x"7C";
END IF;
END BUCLE_INI;
-------------------

------BUCLE_FIN()----
----------------------
FUNCTION BUCLE_FIN(DATO9 : INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT7 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF DATO9 = 1 THEN RETURN '1'&x"7D";
ELSE RETURN '1'&x"7D";
END IF;
END BUCLE_FIN;
-------------------

------LIMPIAR_PANTALLA()----
----------------------
FUNCTION LIMPIAR_PANTALLA(DATO9 : STD_LOGIC)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT10 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF DATO9 = '1' THEN RETURN '1'&x"FE";
ELSE RETURN '1'&x"FD";
END IF;
END LIMPIAR_PANTALLA;
-------------------

------CHAR_ASCII()----
----------------------
FUNCTION CHAR_ASCII(DATO6 : STD_LOGIC_VECTOR(7 DOWNTO 0))RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT4 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
DATAOUT4 := '0'&DATO6;
RETURN DATAOUT4;

END CHAR_ASCII;
-------------------

------CREAR_CHAR()----
----------------------
FUNCTION CREAR_CHAR(DATO11: INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT8 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF 	DATO11 = 1 THEN RETURN '1'&x"7E";
ELSIF DATO11 = 2 THEN RETURN '1'&x"7F";
ELSIF DATO11 = 3 THEN RETURN '1'&x"80";
ELSIF DATO11 = 4 THEN RETURN '1'&x"81";
ELSIF DATO11 = 5 THEN RETURN '1'&x"82";
ELSIF DATO11 = 6 THEN RETURN '1'&x"83";
ELSIF DATO11 = 7 THEN RETURN '1'&x"84";
ELSIF DATO11 = 8 THEN RETURN '1'&x"85";
ELSE RETURN '1'&X"85";
END IF;
END CREAR_CHAR;
-------------------

--------CHAR_CREADO()----
------------------------
FUNCTION CHAR_CREADO(DATO12:INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT9 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF 	DATO12 = 1 THEN RETURN '1'&x"86";
ELSIF DATO12 = 2 THEN RETURN '1'&x"87";
ELSIF DATO12 = 3 THEN RETURN '1'&x"88";
ELSIF DATO12 = 4 THEN RETURN '1'&x"89";
ELSIF DATO12 = 5 THEN RETURN '1'&x"8A";
ELSIF DATO12 = 6 THEN RETURN '1'&x"8B";
ELSIF DATO12 = 7 THEN RETURN '1'&x"8C";
ELSIF DATO12 = 8 THEN RETURN '1'&x"8D";
ELSE  RETURN '1'&x"8D";
END IF;
END CHAR_CREADO;
---------------------

------CODIGO_FIN()----
----------------------
FUNCTION CODIGO_FIN(DATO7 : INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT5 : STD_LOGIC_VECTOR(8 DOWNTO 0);
BEGIN
IF DATO7 = 1 THEN RETURN '1'&x"FF";
ELSE RETURN '1'&x"FF";
END IF;
END CODIGO_FIN;
-------------------
 
end COMANDOS_LCD_REVB;
